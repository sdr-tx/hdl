`include "../../inc/project_defines.v"

module modulator #(
    parameter FOO = 10,
    parameter AM_CLKS_IN_PWM_STEPS = `AM_CLKS_IN_PWM_STEPS,
    parameter AM_PWM_STEPS = `AM_PWM_STEPS
)(
    input clk,
    input rst,
    output pwm
);
    localparam WIDTH = $clog2(FOO);

    /* registers */
    reg [WIDTH-1:0] count;
    wire tc_pwm_step, tc_pwm_symb;
    reg [AM_PWM_STEPS-1:0] shift_register;


    /******** testing signals ********/
    reg [10:0] counter_sine_1k;
    
    /******** testing signals ********/


    // counter to generate ticks at pwm-steps frequency
    counter #(
        .MODULE  (`AM_CLKS_IN_PWM_STEPS)
    ) inst_counter_pwm_steps (
        .clk    (clk),
        .rst    (rst),
        .enable (1'b1),
        .tc     (tc_pwm_step)
    );

    // counter to generate ticks at pwm-symbols frequency
    counter #(
        .MODULE  (AM_PWM_STEPS)
    ) inst_counter_pwm_symb (
        .clk    (clk),
        .rst    (rst),
        .enable (tc_pwm_step),
        .tc     (tc_pwm_symb)
    );

    // shift register to serialize each pwm-symbol
    always @ (posedge clk) begin
        if(rst == 1'b1)begin
            shift_register =0;
            counter_sine_1k <= 0;

        end  else if (tc_pwm_symb == 1'b1) begin
            if(counter_sine_1k == 10'd1000)
                counter_sine_1k = 0;
            else begin
                counter_sine_1k <= counter_sine_1k + 1;

                case(counter_sine_1k)

                10'd0:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd1:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd2:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd3:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd4:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd5:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd6:   shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd7:   shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd8:   shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd9:   shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd10:  shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd11:  shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd12:  shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd13:  shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd14:  shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd15:  shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd16:  shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd17:  shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd18:  shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd19:  shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd20:  shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd21:  shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd22:  shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd23:  shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd24:  shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd25:  shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd26:  shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd27:  shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd28:  shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd29:  shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd30:  shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd31:  shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd32:  shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd33:  shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd34:  shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd35:  shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd36:  shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd37:  shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd38:  shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd39:  shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd40:  shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd41:  shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd42:  shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd43:  shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd44:  shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd45:  shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd46:  shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd47:  shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd48:  shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd49:  shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd50:  shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd51:  shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd52:  shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd53:  shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd54:  shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd55:  shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd56:  shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd57:  shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd58:  shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd59:  shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd60:  shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd61:  shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd62:  shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd63:  shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd64:  shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd65:  shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd66:  shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd67:  shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd68:  shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd69:  shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd70:  shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd71:  shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd72:  shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd73:  shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd74:  shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd75:  shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd76:  shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd77:  shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd78:  shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd79:  shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd80:  shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd81:  shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd82:  shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd83:  shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd84:  shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd85:  shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd86:  shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd87:  shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd88:  shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd89:  shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd90:  shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd91:  shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd92:  shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd93:  shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd94:  shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd95:  shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd96:  shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd97:  shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd98:  shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd99:  shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd100: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd101: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd102: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd103: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd104: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd105: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd106: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd107: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd108: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd109: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd110: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd111: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd112: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd113: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd114: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd115: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd116: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd117: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd118: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd119: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd120: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd121: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd122: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd123: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd124: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd125: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd126: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd127: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd128: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd129: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd130: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd131: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd132: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd133: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd134: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd135: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd136: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd137: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd138: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd139: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd140: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd141: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd142: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd143: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd144: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd145: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd146: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd147: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd148: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd149: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd150: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd151: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd152: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd153: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd154: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd155: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd156: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd157: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd158: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd159: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd160: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd161: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd162: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd163: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd164: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd165: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd166: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd167: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd168: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd169: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd170: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd171: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd172: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd173: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd174: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd175: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd176: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd177: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd178: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd179: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd180: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd181: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd182: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd183: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd184: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd185: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd186: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd187: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd188: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd189: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd190: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd191: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd192: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd193: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd194: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd195: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd196: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd197: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd198: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd199: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd200: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd201: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd202: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd203: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd204: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd205: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd206: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd207: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd208: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd209: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd210: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd211: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd212: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd213: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd214: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd215: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd216: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd217: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd218: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd219: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd220: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd221: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd222: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd223: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd224: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd225: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd226: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd227: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd228: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd229: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd230: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd231: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd232: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd233: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd234: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd235: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd236: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd237: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd238: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd239: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd240: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd241: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd242: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd243: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd244: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd245: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd246: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd247: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd248: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd249: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd250: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd251: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd252: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd253: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd254: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd255: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd256: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd257: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd258: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd259: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd260: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd261: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd262: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd263: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd264: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd265: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd266: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd267: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd268: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd269: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd270: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd271: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd272: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd273: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd274: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd275: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd276: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd277: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd278: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                10'd279: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd280: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd281: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd282: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd283: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd284: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd285: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd286: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd287: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd288: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd289: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd290: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd291: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd292: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd293: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd294: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd295: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd296: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd297: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd298: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd299: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                10'd300: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd301: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd302: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd303: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd304: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd305: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd306: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd307: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd308: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd309: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd310: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd311: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd312: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd313: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                10'd314: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd315: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd316: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd317: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd318: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd319: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd320: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd321: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd322: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd323: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd324: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd325: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                10'd326: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd327: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd328: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd329: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd330: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd331: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd332: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd333: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd334: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd335: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd336: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                10'd337: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd338: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd339: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd340: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd341: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd342: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd343: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd344: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd345: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                10'd346: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd347: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd348: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd349: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd350: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd351: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd352: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd353: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd354: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                10'd355: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd356: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd357: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd358: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd359: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd360: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd361: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd362: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                10'd363: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd364: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd365: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd366: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd367: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd368: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd369: shift_register <= 64'b1111111111111111111111111111111111111111111111111111111000000000;
                10'd370: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd371: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd372: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd373: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd374: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd375: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd376: shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                10'd377: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd378: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd379: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd380: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd381: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd382: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd383: shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                10'd384: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd385: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd386: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd387: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd388: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd389: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd390: shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                10'd391: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd392: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd393: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd394: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd395: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd396: shift_register <= 64'b1111111111111111111111111111111111111111111111111110000000000000;
                10'd397: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd398: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd399: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd400: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd401: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd402: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd403: shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                10'd404: shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd405: shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd406: shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd407: shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd408: shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd409: shift_register <= 64'b1111111111111111111111111111111111111111111111111000000000000000;
                10'd410: shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd411: shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd412: shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd413: shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd414: shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd415: shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                10'd416: shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd417: shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd418: shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd419: shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd420: shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd421: shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                10'd422: shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd423: shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd424: shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd425: shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd426: shift_register <= 64'b1111111111111111111111111111111111111111111111000000000000000000;
                10'd427: shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd428: shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd429: shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd430: shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd431: shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd432: shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                10'd433: shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd434: shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd435: shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd436: shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd437: shift_register <= 64'b1111111111111111111111111111111111111111111100000000000000000000;
                10'd438: shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd439: shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd440: shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd441: shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd442: shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd443: shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                10'd444: shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd445: shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd446: shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd447: shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd448: shift_register <= 64'b1111111111111111111111111111111111111111110000000000000000000000;
                10'd449: shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd450: shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd451: shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd452: shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd453: shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                10'd454: shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd455: shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd456: shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd457: shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd458: shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd459: shift_register <= 64'b1111111111111111111111111111111111111111000000000000000000000000;
                10'd460: shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd461: shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd462: shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd463: shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd464: shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                10'd465: shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd466: shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd467: shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd468: shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd469: shift_register <= 64'b1111111111111111111111111111111111111100000000000000000000000000;
                10'd470: shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd471: shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd472: shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd473: shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd474: shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                10'd475: shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd476: shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd477: shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd478: shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd479: shift_register <= 64'b1111111111111111111111111111111111110000000000000000000000000000;
                10'd480: shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd481: shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd482: shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd483: shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd484: shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                10'd485: shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd486: shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd487: shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd488: shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd489: shift_register <= 64'b1111111111111111111111111111111111000000000000000000000000000000;
                10'd490: shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd491: shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd492: shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd493: shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd494: shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                10'd495: shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd496: shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd497: shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd498: shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd499: shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd500: shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                10'd501: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd502: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd503: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd504: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd505: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd506: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd507: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd508: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd509: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd510: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd511: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd512: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd513: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd514: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd515: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd516: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd517: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd518: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd519: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd520: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd521: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd522: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd523: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd524: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd525: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd526: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd527: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd528: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd529: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd530: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd531: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd532: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd533: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd534: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd535: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd536: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd537: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd538: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd539: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd540: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd541: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd542: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd543: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd544: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd545: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd546: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd547: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd548: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd549: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd550: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd551: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd552: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd553: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd554: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd555: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd556: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd557: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd558: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd559: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd560: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd561: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd562: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd563: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd564: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd565: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd566: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd567: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd568: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd569: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd570: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd571: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd572: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd573: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd574: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd575: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd576: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd577: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd578: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd579: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd580: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd581: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd582: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd583: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd584: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd585: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd586: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd587: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd588: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd589: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd590: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd591: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd592: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd593: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd594: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd595: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd596: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd597: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd598: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd599: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd600: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd601: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd602: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd603: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd604: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd605: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd606: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd607: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd608: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd609: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd610: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd611: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd612: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd613: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd614: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd615: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd616: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd617: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd618: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd619: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd620: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd621: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd622: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd623: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd624: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd625: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd626: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd627: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd628: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd629: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd630: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd631: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd632: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd633: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd634: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd635: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd636: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd637: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd638: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd639: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd640: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd641: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd642: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd643: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd644: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd645: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd646: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd647: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd648: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd649: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd650: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd651: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd652: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd653: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd654: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd655: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd656: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd657: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd658: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd659: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd660: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd661: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd662: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd663: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd664: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd665: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd666: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd667: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd668: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd669: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd670: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd671: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd672: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd673: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd674: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd675: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd676: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd677: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd678: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd679: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd680: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd681: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd682: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd683: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd684: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd685: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd686: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd687: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd688: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd689: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd690: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd691: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd692: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd693: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd694: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd695: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd696: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd697: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd698: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd699: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd700: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd701: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd702: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd703: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd704: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd705: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd706: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd707: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd708: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd709: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd710: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd711: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd712: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd713: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd714: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd715: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd716: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd717: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd718: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd719: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd720: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd721: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd722: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd723: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd724: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd725: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd726: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd727: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd728: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd729: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd730: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd731: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd732: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd733: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd734: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd735: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd736: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd737: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd738: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd739: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd740: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd741: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd742: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd743: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd744: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd745: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd746: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd747: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd748: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd749: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd750: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd751: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd752: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd753: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd754: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd755: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd756: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd757: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd758: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd759: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd760: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd761: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd762: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd763: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd764: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd765: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd766: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd767: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd768: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd769: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd770: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd771: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd772: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd773: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd774: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd775: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd776: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd777: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd778: shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                10'd779: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd780: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd781: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd782: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd783: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd784: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd785: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd786: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd787: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd788: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd789: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd790: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd791: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd792: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd793: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd794: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd795: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd796: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd797: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd798: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd799: shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                10'd800: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd801: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd802: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd803: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd804: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd805: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd806: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd807: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd808: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd809: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd810: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd811: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd812: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd813: shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                10'd814: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd815: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd816: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd817: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd818: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd819: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd820: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd821: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd822: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd823: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd824: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd825: shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                10'd826: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd827: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd828: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd829: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd830: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd831: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd832: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd833: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd834: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd835: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd836: shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                10'd837: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd838: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd839: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd840: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd841: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd842: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd843: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd844: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd845: shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                10'd846: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd847: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd848: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd849: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd850: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd851: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd852: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd853: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd854: shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                10'd855: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd856: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd857: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd858: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd859: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd860: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd861: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd862: shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                10'd863: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd864: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd865: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd866: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd867: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd868: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd869: shift_register <= 64'b1111111100000000000000000000000000000000000000000000000000000000;
                10'd870: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd871: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd872: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd873: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd874: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd875: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd876: shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                10'd877: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd878: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd879: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd880: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd881: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd882: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd883: shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                10'd884: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd885: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd886: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd887: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd888: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd889: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd890: shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                10'd891: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd892: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd893: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd894: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd895: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd896: shift_register <= 64'b1111111111110000000000000000000000000000000000000000000000000000;
                10'd897: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd898: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd899: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd900: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd901: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd902: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd903: shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                10'd904: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd905: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd906: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd907: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd908: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd909: shift_register <= 64'b1111111111111100000000000000000000000000000000000000000000000000;
                10'd910: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd911: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd912: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd913: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd914: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd915: shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                10'd916: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd917: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd918: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd919: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd920: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd921: shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                10'd922: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd923: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd924: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd925: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd926: shift_register <= 64'b1111111111111111100000000000000000000000000000000000000000000000;
                10'd927: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd928: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd929: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd930: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd931: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd932: shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                10'd933: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd934: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd935: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd936: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd937: shift_register <= 64'b1111111111111111111000000000000000000000000000000000000000000000;
                10'd938: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd939: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd940: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd941: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd942: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd943: shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                10'd944: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd945: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd946: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd947: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd948: shift_register <= 64'b1111111111111111111110000000000000000000000000000000000000000000;
                10'd949: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd950: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd951: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd952: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd953: shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                10'd954: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd955: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd956: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd957: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd958: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd959: shift_register <= 64'b1111111111111111111111100000000000000000000000000000000000000000;
                10'd960: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd961: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd962: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd963: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd964: shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                10'd965: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd966: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd967: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd968: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd969: shift_register <= 64'b1111111111111111111111111000000000000000000000000000000000000000;
                10'd970: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd971: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd972: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd973: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd974: shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                10'd975: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd976: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd977: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd978: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd979: shift_register <= 64'b1111111111111111111111111110000000000000000000000000000000000000;
                10'd980: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd981: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd982: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd983: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd984: shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                10'd985: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd986: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd987: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd988: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd989: shift_register <= 64'b1111111111111111111111111111100000000000000000000000000000000000;
                10'd990: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd991: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd992: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd993: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd994: shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                10'd995: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd996: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd997: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd998: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                10'd999: shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
        
                default:
                    shift_register <= 64'd0;
    
                endcase
            end

        end else if (tc_pwm_step == 1'b1)
            shift_register <= {shift_register[AM_PWM_STEPS-2:0],shift_register[AM_PWM_STEPS-1]};

    end

    // output assignment
    assign pwm = shift_register[AM_PWM_STEPS-1];


endmodule


