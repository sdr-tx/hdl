`include "../../inc/project_defines.v"

module modulator #(
    parameter FOO = 10,
    parameter AM_CLKS_IN_PWM_STEPS = `AM_CLKS_IN_PWM_STEPS,
    parameter AM_PWM_STEPS = `AM_PWM_STEPS
)(
    input clk,
    input rst,
    output pwm
);
    localparam WIDTH = $clog2(FOO);

    /* registers */
    reg [WIDTH-1:0] count;
    wire tc_pwm_step, tc_pwm_symb;
    reg [AM_PWM_STEPS-1:0] shift_register;


    /******** testing signals ********/
/*    localparam [6:0] sine_10
    {
32'h428a2f98,32'h71374491,32'hb5c0fbcf,32'he9b5dba5,32'h3956c25b,32'h59f111f1,32'h923f82a4,32'hab1c5ed5,
32'hd807aa98,32'h12835b01,32'h243185be,32'h550c7dc3,32'h72be5d74,32'h80deb1fe,32'h9bdc06a7,32'hc19bf174,
32'he49b69c1,32'hefbe4786,32'h0fc19dc6,32'h240ca1cc,32'h2de92c6f,32'h4a7484aa,32'h5cb0a9dc,32'h76f988da,
32'h983e5152,32'ha831c66d,32'hb00327c8,32'hbf597fc7,32'hc6e00bf3,32'hd5a79147,32'h06ca6351,32'h14292967,
32'h27b70a85,32'h2e1b2138,32'h4d2c6dfc,32'h53380d13,32'h650a7354,32'h766a0abb,32'h81c2c92e,32'h92722c85,
32'ha2bfe8a1,32'ha81a664b,32'hc24b8b70,32'hc76c51a3,32'hd192e819,32'hd6990624,32'hf40e3585,32'h106aa070,
32'h19a4c116,32'h1e376c08,32'h2748774c,32'h34b0bcb5,32'h391c0cb3,32'h4ed8aa4a,32'h5b9cca4f,32'h682e6ff3,
32'h748f82ee,32'h78a5636f,32'h84c87814,32'h8cc70208,32'h90befffa,32'ha4506ceb,32'hbef9a3f7,32'hc67178f2
};*/
    reg [6:0] counter_sine_10k;
    /******** testing signals ********/


    // counter to generate ticks at pwm-steps frequency
    counter #(
        .MODULE  (`AM_CLKS_IN_PWM_STEPS)
    ) inst_counter_pwm_steps (
        .clk    (clk),
        .rst    (rst),
        .enable (1'b1),
        .tc     (tc_pwm_step)
    );

    // counter to generate ticks at pwm-symbols frequency
    counter #(
        .MODULE  (AM_PWM_STEPS)
    ) inst_counter_pwm_symb (
        .clk    (clk),
        .rst    (rst),
        .enable (tc_pwm_step),
        .tc     (tc_pwm_symb)
    );

    // shift register to serialize each pwm-symbol
    always @ (posedge clk) begin
        if(rst == 1'b1)begin
            shift_register <= `AM_PWM_STEPS'd0;
            counter_sine_10k <= 0;
        end
        else if (tc_pwm_symb == 1'b1) begin
            if(counter_sine_10k == 7'd100)
                counter_sine_10k = 7'd0;
            else begin
                counter_sine_10k <= counter_sine_10k + 1;
                case(counter_sine_10k)
                    // 0 - 10
                    7'd0:   shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                    7'd1:   shift_register <= 64'b1111111111111111111111111111111100000000000000000000000000000000;
                    7'd2:   shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                    7'd3:   shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                    7'd4:   shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                    7'd5:   shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                    7'd6:   shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                    7'd7:   shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                    7'd8:   shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                    7'd9:   shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                    7'd10:   shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                    7'd11:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                    7'd12:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                    7'd13:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                    7'd14:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                    7'd15:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                    7'd16:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                    7'd17:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                    7'd18:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                    7'd19:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                    7'd20:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                    7'd21:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                    7'd22:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                    7'd23:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    7'd24:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    7'd25:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    7'd26:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    7'd27:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    7'd28:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                    7'd29:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111100;
                    7'd30:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                    7'd31:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111111000;
                    7'd32:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111110000;
                    7'd33:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111100000;
                    7'd34:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111111000000;
                    7'd35:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111110000000;
                    7'd36:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111111100000000;
                    7'd37:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111110000000000;
                    7'd38:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111100000000000;
                    7'd39:   shift_register <= 64'b1111111111111111111111111111111111111111111111111111000000000000;
                    7'd40:   shift_register <= 64'b1111111111111111111111111111111111111111111111111100000000000000;
                    7'd41:   shift_register <= 64'b1111111111111111111111111111111111111111111111110000000000000000;
                    7'd42:   shift_register <= 64'b1111111111111111111111111111111111111111111111100000000000000000;
                    7'd43:   shift_register <= 64'b1111111111111111111111111111111111111111111110000000000000000000;
                    7'd44:   shift_register <= 64'b1111111111111111111111111111111111111111111000000000000000000000;
                    7'd45:   shift_register <= 64'b1111111111111111111111111111111111111111100000000000000000000000;
                    7'd46:   shift_register <= 64'b1111111111111111111111111111111111111110000000000000000000000000;
                    7'd47:   shift_register <= 64'b1111111111111111111111111111111111111000000000000000000000000000;
                    7'd48:   shift_register <= 64'b1111111111111111111111111111111111100000000000000000000000000000;
                    7'd49:   shift_register <= 64'b1111111111111111111111111111111110000000000000000000000000000000;
                    7'd50:   shift_register <= 64'b1111111111111111111111111111111000000000000000000000000000000000;
                    7'd51:   shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;
                    7'd52:   shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                    7'd53:   shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                    7'd54:   shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                    7'd55:   shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                    7'd56:   shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                    7'd57:   shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                    7'd58:   shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                    7'd59:   shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                    7'd60:   shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                    7'd61:   shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                    7'd62:   shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                    7'd63:   shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                    7'd64:   shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                    7'd65:   shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                    7'd66:   shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                    7'd67:   shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                    7'd68:   shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                    7'd69:   shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                    7'd70:   shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                    7'd71:   shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                    7'd72:   shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                    7'd73:   shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7'd74:   shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7'd75:   shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7'd76:   shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7'd77:   shift_register <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7'd78:   shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                    7'd79:   shift_register <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
                    7'd80:   shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                    7'd81:   shift_register <= 64'b1100000000000000000000000000000000000000000000000000000000000000;
                    7'd82:   shift_register <= 64'b1110000000000000000000000000000000000000000000000000000000000000;
                    7'd83:   shift_register <= 64'b1111000000000000000000000000000000000000000000000000000000000000;
                    7'd84:   shift_register <= 64'b1111100000000000000000000000000000000000000000000000000000000000;
                    7'd85:   shift_register <= 64'b1111110000000000000000000000000000000000000000000000000000000000;
                    7'd86:   shift_register <= 64'b1111111000000000000000000000000000000000000000000000000000000000;
                    7'd87:   shift_register <= 64'b1111111110000000000000000000000000000000000000000000000000000000;
                    7'd88:   shift_register <= 64'b1111111111000000000000000000000000000000000000000000000000000000;
                    7'd89:   shift_register <= 64'b1111111111100000000000000000000000000000000000000000000000000000;
                    7'd90:   shift_register <= 64'b1111111111111000000000000000000000000000000000000000000000000000;
                    7'd91:   shift_register <= 64'b1111111111111110000000000000000000000000000000000000000000000000;
                    7'd92:   shift_register <= 64'b1111111111111111000000000000000000000000000000000000000000000000;
                    7'd93:   shift_register <= 64'b1111111111111111110000000000000000000000000000000000000000000000;
                    7'd94:   shift_register <= 64'b1111111111111111111100000000000000000000000000000000000000000000;
                    7'd95:   shift_register <= 64'b1111111111111111111111000000000000000000000000000000000000000000;
                    7'd96:   shift_register <= 64'b1111111111111111111111110000000000000000000000000000000000000000;
                    7'd97:   shift_register <= 64'b1111111111111111111111111100000000000000000000000000000000000000;
                    7'd98:   shift_register <= 64'b1111111111111111111111111111000000000000000000000000000000000000;
                    7'd99:   shift_register <= 64'b1111111111111111111111111111110000000000000000000000000000000000;

                    default:
                        shift_register <= 64'd0;                    
                endcase
            end
        end else if (tc_pwm_step == 1'b1)
            shift_register <= {shift_register[AM_PWM_STEPS-2:0],shift_register[AM_PWM_STEPS-1]};
    end

    // output assignment
    assign pwm = shift_register[AM_PWM_STEPS-1];

endmodule


